module constant #(parameter VALUE = 4) (
    output [31:0] out
);

assign out = VALUE;

endmodule
